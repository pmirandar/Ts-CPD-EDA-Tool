- op-amp, main
* 
*
.include param.cir
*.include opamp-main.cir
* opamp desciption
* power supplies
VDD 4 0 DC +5V
Vss 5 0 DC -5V
*Vc1 2 0 DC 1.2V
*Vc2 5 0 DC 1.2V
* differential-mode signal level
*Vd 21 0 DC 0V
Vd 101 0 sin(0 0.1 100000000) ac 1.0V dc 0.0
*Vd 21 0 dc 0.0 ac 1 0
*+ distof1 1 0
*+ distof2 1 0
*+ sin(0 0.1V 100000000 0 0)
*vin 2 5 sin(0 0.1 20000000) ac 1.0V dc 0.0
* to DC sweep the input common-mode level, offset diff-input by +220uV
*Vd 21 0 DC +220.0uV
Rd 101 0 1
EV1 2 100 101 0 +0.5
EV2 1 100 101 0 -0.5
*EV1 2 100 101 0 +1.0
*EV2 1 100 101 0 -1.0
* common-mode signal level
Vcm 100 0 DC 0V
* front-end stage
M2 6 9 4 4 CMOSP L=1.6u W={w2}
M3 7 1 6 4 CMOSP L=1.6u W={w3}
M4 8 2 6 4 CMOSP L=1.6u W={w4}
M5 7 7 5 5 CMOSN L=1.6u W={w5}
M6 8 7 5 5 CMOSN L=1.6u W={w6}
* 2nd gain stage
M7 3 9 4 4 CMOSP L=1.6u W={w7}
M8 3 8 5 5 CMOSN L=1.6u W={w8}
* current source biasing stage
M1 9 9 4 4 CMOSP L=1.6u W={w1}
Iref 9 5 dc 20uA
* compensation network
Rc 10 3 {Rc}
Cc 8 10 {CAPc}
* load for the op-amp
CL 3 0 1.0pF
.model CMOSN  nmos Version=3.2.2
+ level=8
+ Tnom=27.0
+ nch= 1.024685E+17  tox=1.00000E-08 xj=1.00000E-07
+ lint= 3.75860E-08 wint=-2.02101528644562E-07
+ vth0= .6094574   k1= .5341038  k2= 1.703463E-03  k3=-17.24589
+ dvt0= .1767506  dvt1= .5109418  dvt2=-0.05
+ nlx= 9.979638E-08  w0=1e-6
+ k3b= 4.139039
+ vsat= 97662.05  ua=-1.748481E-09  ub= 3.178541E-18  uc=1.3623e-10
+ rdsw= 298.873  u0= 307.2991 prwb=-2.24e-4
+ a0= .4976366
+ keta=-2.195445E-02  a1= .0332883  a2= .9
+ voff=-9.623903E-02  nFactor= .8408191  cit= 3.994609E-04
+ cdsc= 1.130797E-04
+ cdscb=2.4e-5
+ eta0= .0145072  etab=-3.870303E-03
+ dsub= .4116711
+ pclm= 1.813153  pdiblc1= 2.003703E-02  pdiblc2= .00129051 pdiblcb=-1.034e-3
+ drout= .4380235  pscbe1= 5.752058E+08  pscbe2= 7.510319E-05
+ pvag= .6370527 prt=68.7 ngate=1.e20 alpha0=1.e-7 beta0=28.4
+ prwg=-0.001 ags=1.2
+ dvt0w=0.58 dvt1w=5.3e6 dvt2w=-0.0032
+ kt1=-.3  kt2=-.03
+ at= 33000
+ ute=-1.5
+ ua1= 4.31E-09  ub1= 7.61E-18  uc1=-2.378e-10
+ kt1l=1e-8
+ wr=1 b0=1e-7 b1=1e-7 dwg=5e-8 dwb=2e-8 delta=0.015
+ cgdl=1e-10 cgsl=1e-10 cgbo=1e-10 xpart=0.0
+ cgdo=0.4e-9 cgso=0.4e-9
+ clc=0.1e-6
+ cle=0.6
+ ckappa=0.6

.model CMOSP  pmos Version=3.2.2
+ level=8
+ Tnom=27.0
+ nch= 5.73068E+16  tox=1.00000E-08 xj=1.00000E-07
+ lint= 8.195860E-08 wint=-1.821562E-07
+ vth0= -.86094574   k1= .341038  k2= 2.703463E-02  k3=12.24589
+ dvt0= .767506  dvt1= .65109418  dvt2=-0.145
+ nlx= 1.979638E-07  w0=1.1e-6
+ k3b= -2.4139039
+ vsat= 60362.05  ua=1.348481E-09  ub= 3.178541E-19  uc=1.1623e-10
+ rdsw= 498.873  u0= 137.2991 prwb=-1.2e-5
+ a0= .3276366
+ keta=-1.8195445E-02  a1= .0232883  a2= .9
+ voff=-6.623903E-02  nFactor= 1.0408191  cit= 4.994609E-04
+ cdsc= 1.030797E-3
+ cdscb=2.84e-4
+ eta0= .0245072  etab=-1.570303E-03
+ dsub= .24116711
+ pclm= 2.6813153  pdiblc1= 4.003703E-02  pdiblc2= .00329051 pdiblcb=-2.e-4
+ drout= .1380235  pscbe1= 0  pscbe2=1.e-28
+ pvag= -.16370527
+ prwg=-0.001 ags=1.2
+ dvt0w=0.58 dvt1w=5.3e6 dvt2w=-0.0032
+ kt1=-.3  kt2=-.03 prt=76.4
+ at= 33000
+ ute=-1.5
+ ua1= 4.31E-09  ub1= 7.61E-18  uc1=-2.378e-10
+ kt1l=0
+ wr=1 b0=1e-7 b1=1e-7 dwg=5e-8 dwb=2e-8 delta=0.015
+ cgdl=1e-10 cgsl=1e-10 cgbo=1e-10 xpart=0.0
+ cgdo=0.4e-9 cgso=0.4e-9
+ clc=0.1e-6
+ cle=0.6
+ ckappa=0.6
*
*** Analysis Requests **
.control
set units=degrees
 OP
** .TF V(13) Vd
*** AC
 tf V(3) Vd
 AC dec 1000 1 80MEGHZ 
* .acphace 0
* Output Requests **
**plot  vdb(3) vp(3)
wrdata ngspice vdb(3) vp(3)
show m6 > m6.data
.endc
.end
