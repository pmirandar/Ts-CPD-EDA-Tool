- op-amp
* 
*
** Circuit Description **
.include SimInOut/param.cir
.options badmos3
.include SimIn/modeloBSIM.cir
.include SimIn/opamp-main-2.cir
*.include SimIn/power-supplies.cir
* power supplies
*vdi={vd}
*vsi={vs}
VDD 4 0 DC +2.5V 
*Vss 5 0 DC 0V
Vss 5 0 DC -2.5V
* differential-mode signal level
*Vd 21 0 DC 0V
Vd 101 0 sin(0 0.1 100000000) ac 1.0V dc +0.8uV
*Vd 21 0 dc 0.0 ac 1 0
*+ distof1 1 0
*+ distof2 1 0
*+ sin(0 0.1V 100000000 0 0)
*vin 2 5 sin(0 0.1 20000000) ac 1.0V dc 0.0
* to DC sweep the input common-mode level, offset diff-input by +220uV
*Vd 21 0 DC +220.0uV
Rd 101 0 1
EV1 2 100 101 0 +0.5
EV2 1 100 101 0 -0.5
* common-mode signal level
Vcm 100 0 DC 0V
*** Analysis Requests **
.control
set units=degrees
 OP
*** AC
 tf V(3) Vd
 AC dec 1000 1 100MEGHZ 
* Output Requests **
wrdata SimInOut/ngspice vdb(3) unwrap(vp(3))
.endc
.end
