.param w1=2e-06 w2=2e-06 w3=2.2853e-06 w4=2.2853e-06 w5=4.6698e-06 w6=4.6698e-06 w7=4.6629e-05 w8=9.9852e-06 CL=1.1996e-11 CAPc=3.1717e-12 l1=2e-06 l2=2e-06 l3=2e-06 l4=2e-06 l5=2e-06 l6=2e-06 l7=2e-06 l8=2e-06 Iref=3.685e-05
