.param w1=1.2674e-05 w2=1.2674e-05 w3=1.8644e-05 w4=1.8644e-05 w5=7.2041e-06 w6=7.2041e-06 w7=3.9366e-05 w8=3.4629e-05 CL=7.4751e-12 CAPc=1.3411e-11 l1=8e-07 l2=8e-07 l3=8e-07 l4=8e-07 l5=8e-07 l6=8e-07 l7=8e-07 l8=8e-07 Iref=4.0383e-05
