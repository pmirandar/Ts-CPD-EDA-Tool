- op-amp
* for calculation of negative Power Supply Rejection Ratio (PSRR-) 
*
.include SimInOut/param.cir
.options badmos3
*.include modelos.mod
.include SimIn/modeloBSIM.cir
.include SimIn/opamp-main-2.cir
* power supplies
VDD 4 0 DC +2.5V
Vss 25 0 DC -2.5V
* Other external connections
Vshort 1 3 0
*Vshort 2 0 0
*Vgnd 2 0 +20 uV
Vgnd 2 0 0
*Vgnd 1 3 0
*Vd 5 25 sin(0 0.1 100000000) ac -1.0V dc 0.8e-6
Vd 5 25 sin(0 0.1 100000000) ac -1.0V dc 0
.control
set units=degrees
OP
*** Analysis Requests **
 AC dec 1000 1 100MEGHZ 
*
* Output Requests **
*plot v(3)
wrdata SimInOut/psrr- v(3)
.endc
.end
