 opamp
* for calculation of slew rate 
*
.include SimInOut/param.cir
*.include modelos.mod
.include SimIn/modeloBSIM.cir
.include SimIn/opamp-main-2.cir
* power supplies
VDD 4 0 DC +2.5V
Vss 5 0 DC -2.5V
Vd 2 0 PWL(0, 0V 1ns,+2.0V 5000ns,+2.0V 5001ns,0V 0.5s, 0V )
* nodo 1 es negativo (-)
Vshort 1 3 0
*                                                            
*** Analysis Requests **
.control
*OP
*tran 100ns 5us
tran 100ns 10us
* Output Requests **
*plot v(2) v(3)
wrdata SimInOut/slewrate v(2) v(3)
.endc
.end
