.param w1=7.1894e-05 w2=7.1894e-05 w3=6.5892e-05 w4=1.3276e-05 w5=1.3276e-05 w6=2.5197e-05 w7=2.5197e-05 w8=8.2574e-05 w9=8.2574e-05 w10=8.2574e-05 w11=8.2574e-05 w12=0.00011166 w13=2.5197e-05 w14=1.3276e-05 w15=1.6933e-05 CL=1e-11 l1=1.25e-06 l2=1.25e-06 l3=1.25e-06 l4=1.25e-06 l5=1.25e-06 l6=1.25e-06 l7=1.25e-06 l8=1.25e-06 l9=1.25e-06 l10=1.25e-06 l11=1.25e-06 l12=1.25e-06 l13=1.25e-06 l14=1.25e-06 l15=1.25e-06 Iref=6.3285e-05 Re1=1659.3458 Re2=1659.3458
