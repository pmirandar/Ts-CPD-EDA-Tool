.param w1=5.4745e-06 w2=7.0241e-05 w3=5.1035e-05 w4=5.1035e-05 w5=4.2696e-06 w6=4.2696e-06 CL=8.3036e-12 l1=1.4e-06 l2=1.4e-06 l3=3.5e-06 l4=3.5e-06 l5=3.5e-06 l6=3.5e-06 Iref=6.7009e-05
