.param w1=0.00019145 w2=1.4041e-05 w3=3.4922e-05 w4=3.4922e-05 w5=2.2336e-05 w6=2.2336e-05 CL=1.3237e-11 l1=1.4e-06 l2=1.4e-06 l3=3.5e-06 l4=3.5e-06 l5=3.5e-06 l6=3.5e-06 Iref=2.2341e-05
