.param vd=2.5 vs=-2.5
