- op-amp
*
** Circuit Description **
.include SimInOut/param.cir
.options badmos3
*.include modelos.mod
.include SimIn/modeloBSIM.cir
.include SimIn/opamp-main-2.cir
* power supplies
VDD 24 0 DC +2.5V
Vss 5 0 DC -2.5V
* Other external connections
Vshort 1 3 0
Vgnd 2 0 0 
*Vd 4 24 sin(0 0.1 10000000) ac 1.0V dc -0.8e-6
Vd 4 24 sin(0 0.1 10000000) ac 1.0V dc 0
.control
set units=degrees
OP
*** Analysis Requests **
* tf V(3) Vd
 AC dec 1000 1 100MEGHZ
* Output Requests **
*plot vdb(3)
wrdata SimInOut/psrr+ v(3)
.endc
.end
